.title KiCad schematic
.include "/home/maykol/Documentos/spice/2SA1943.lib"
.include "/home/maykol/Documentos/spice/2SC5200.mod"
.include "/home/maykol/Documentos/spice/2n5401.lib"
.include "/home/maykol/Documentos/spice/2n5551.lib"
.include "/home/maykol/Documentos/spice/Standard_Rectifiers.lib"
.include "/home/maykol/Documentos/spice/transistores_2.lib"
.save all
.probe alli

**comienzo de las pruebas
*.op
.tran 10u 5m 1m
.measure tran Vo_RMS RMS v(/voq103) from=2m to=4m
.measure tran Io_RMS RMS i(R102) from=2m to=4m
.measure tran ir105_RMS RMS i(r105) from=2m to=4m
.measure tran ir104_RMS RMS i(r104) from=2m to=4m
.control
fourier 1k v(/voq103)
gnuplot Vo v(/voq103) v(/v4i)
+ xycontour
+ title 'Voltaje de salida Vs Voltaje de entrada'
+ xlabel 'Tiempo (S)'
+ ylabel 'Voltaje (V)'
.endc

**Fin de las pruebas
V1 +50V GND DC 50 
V2 GND -50V DC 50 
R9 +50V /VE2 150
Q2 /VC2 /VB2 /VE2 2N5401
Q5 Net-_Q4-B_ Net-_Q4-B_ Net-_Q5-E_ 2N5551
R10 Net-_Q4-E_ -50V 68
Q4 Net-_Q4-C_ Net-_Q4-B_ Net-_Q4-E_ 2N5551
R15 Net-_Q5-E_ -50V 68
Q8 Net-_Q4-B_ Net-_Q8-B_ Net-_Q8-E_ 2N5401
R18 /VC2 Net-_Q7-E_ 100
Q7 Net-_Q4-C_ Net-_Q7-B_ Net-_Q7-E_ 2N5401
R11 /VC2 Net-_Q8-E_ 100
C8 -50V GND 100n
C102 Net-_Q7-B_ /v4i 3.3u
V4 /v4i GND DC 0 SIN( 0 2 1k 0 0 0 2 ) AC 2 
R22 Net-_Q7-B_ GND 10k
R14 /VE2 Net-_Q3-B_ 1k
R13 /VB2 /gndv 10k
Q3 /VB2 Net-_Q3-B_ +50V 2N5401
C3 +50V /gndv 10u
R12 /gndv GND 12k
R101 +50V Net-_Q102-E_ 100
Q102 /vdt /VB2 Net-_Q102-E_ 2N5401
Q112 /vdt Net-_Q112-B_ /vdb 2N5551
R115 /vdt Net-_Q112-B_ 1.2k
Q103 +50V /vdt Net-_Q10-B_ 2SD669
R21 Net-_Q9-E_ -50V 22
Q9 /vdb Net-_Q4-C_ Net-_Q9-E_ 2N5551
Q104 -50V /vdb Net-_Q101-B_ 2SB649
R20 Net-_C6-Pad1_ Net-_Q8-B_ 1k
C6 Net-_C6-Pad1_ GND 220u
C5 Net-_Q4-C_ /vdb 300p
R19 Net-_Q8-B_ Net-_C7-Pad1_ 220
R23 Net-_Q8-B_ /voq103 18k
C7 Net-_C7-Pad1_ /voq103 100p
R103 /voq103 Net-_Q101-B_ 33
R116 Net-_Q112-B_ /vdb 330
XQ101 -50V Net-_Q101-B_ Net-_Q101-E_ 2SA1943
R109 /voq103 Net-_Q107-E_ 0.33
R108 Net-_Q106-E_ /voq103 0.33
XQ107 -50V Net-_Q101-B_ Net-_Q107-E_ 2SA1943
Q106 +50V Net-_Q10-B_ Net-_Q106-E_ 2SC5200
R102 /voq103 GND 8
R106 /voq103 Net-_Q101-E_ 0.33
Q10 +50V Net-_Q10-B_ Net-_Q10-E_ 2SC5200
R105 Net-_Q10-E_ /voq103 0.33
R104 Net-_Q10-B_ /voq103 33
.end
